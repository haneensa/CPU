----------------------------------------------------------------------------------
-- Engineer: 
-- Create Date:    13:34:01 12/13/2014 
-- Module Name:    ALU - Behavioral 
-- Description: 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ALU is
end ALU;

architecture Behavioral of ALU is

begin


end Behavioral;

