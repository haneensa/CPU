----------------------------------------------------------------------------------
-- Engineer: 
-- Create Date:    13:34:43 12/13/2014 
-- Module Name:    control_unit - Behavioral 
-- Description: 


----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity control_unit is
end control_unit;

architecture Behavioral of control_unit is

begin


end Behavioral;

