---------------------------------------------------------------------------------- 
-- Engineer: 
-- Create Date:    13:32:21 12/13/2014 
-- Module Name:    instruction_register - Behavioral 
-- Description: 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity instruction_register is
end instruction_register;

architecture Behavioral of instruction_register is

begin


end Behavioral;

