----------------------------------------------------------------------------------
-- Engineer: 
-- Create Date:    13:39:20 12/13/2014 
-- Module Name:    memory_data_register - Behavioral 
-- Description: 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity memory_data_register is
end memory_data_register;

architecture Behavioral of memory_data_register is

begin


end Behavioral;

