----------------------------------------------------------------------------------
-- Engineer: 
-- Create Date:    13:38:42 12/13/2014  
-- Module Name:    memory_address_register - Behavioral 
-- Description: 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity memory_address_register is
end memory_address_register;

architecture Behavioral of memory_address_register is

begin


end Behavioral;

