----------------------------------------------------------------------------------
-- Engineer: 
-- Create Date:    18:36:24 12/15/2014 
-- Module Name:    instruction_decoder - Behavioral 
-- Project Name: 
-- Description: take the instruction from the IR and decode the instruction then sends the 
-- relevent data to ALU or control unit or Registers
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity instruction_decoder is
end instruction_decoder;

architecture Behavioral of instruction_decoder is

begin


end Behavioral;

